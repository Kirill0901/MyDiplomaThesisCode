﻿        None            = 0,    ///< Пустая операция
        PushConst       = 1,    ///< Оператор выкладывания константы на стек
        Assign          = 2,    ///< Оператор присваивания
        Equal           = 3,   ///< Логическое равенство
        NotEqual        = 4,   ///< Логическое неравенство
        Less            = 5,   ///< Логическое меньше
        LessOrEqual     = 6,   ///< Логическое меньше или равно
        More            = 7,   ///< Логическое больше
        MoreOrEqual     = 8,   ///< Логическое больше или равно
